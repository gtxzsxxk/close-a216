module cpu_top(
    input CLK
);

endmodule